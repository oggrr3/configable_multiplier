module ev_generator (
    input   [7:0]   multiplicand_i      ,
    input   [7:0]   multiplier_i        ,
    intput          enable_i            ,
    ouput   [15:0]
);

endmodule